`default_nettype none

module Template
(
  input  logic        clk, reset_n,
  input  logic [11:0] A,
  input  logic        update,
  output logic [11:0] S
);

endmodule: Template