// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: history_reg.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 12.1 Build 177 11/07/2012 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2012 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module history_reg (
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps100x,
	taps101x,
	taps102x,
	taps103x,
	taps104x,
	taps105x,
	taps106x,
	taps107x,
	taps108x,
	taps109x,
	taps10x,
	taps110x,
	taps111x,
	taps112x,
	taps113x,
	taps114x,
	taps115x,
	taps116x,
	taps117x,
	taps118x,
	taps119x,
	taps11x,
	taps120x,
	taps121x,
	taps122x,
	taps123x,
	taps124x,
	taps125x,
	taps126x,
	taps127x,
	taps12x,
	taps13x,
	taps14x,
	taps15x,
	taps16x,
	taps17x,
	taps18x,
	taps19x,
	taps1x,
	taps20x,
	taps21x,
	taps22x,
	taps23x,
	taps24x,
	taps25x,
	taps26x,
	taps27x,
	taps28x,
	taps29x,
	taps2x,
	taps30x,
	taps31x,
	taps32x,
	taps33x,
	taps34x,
	taps35x,
	taps36x,
	taps37x,
	taps38x,
	taps39x,
	taps3x,
	taps40x,
	taps41x,
	taps42x,
	taps43x,
	taps44x,
	taps45x,
	taps46x,
	taps47x,
	taps48x,
	taps49x,
	taps4x,
	taps50x,
	taps51x,
	taps52x,
	taps53x,
	taps54x,
	taps55x,
	taps56x,
	taps57x,
	taps58x,
	taps59x,
	taps5x,
	taps60x,
	taps61x,
	taps62x,
	taps63x,
	taps64x,
	taps65x,
	taps66x,
	taps67x,
	taps68x,
	taps69x,
	taps6x,
	taps70x,
	taps71x,
	taps72x,
	taps73x,
	taps74x,
	taps75x,
	taps76x,
	taps77x,
	taps78x,
	taps79x,
	taps7x,
	taps80x,
	taps81x,
	taps82x,
	taps83x,
	taps84x,
	taps85x,
	taps86x,
	taps87x,
	taps88x,
	taps89x,
	taps8x,
	taps90x,
	taps91x,
	taps92x,
	taps93x,
	taps94x,
	taps95x,
	taps96x,
	taps97x,
	taps98x,
	taps99x,
	taps9x);

	input	  clock;
	input	[11:0]  shiftin;
	output	[11:0]  shiftout;
	output	[11:0]  taps0x;
	output	[11:0]  taps100x;
	output	[11:0]  taps101x;
	output	[11:0]  taps102x;
	output	[11:0]  taps103x;
	output	[11:0]  taps104x;
	output	[11:0]  taps105x;
	output	[11:0]  taps106x;
	output	[11:0]  taps107x;
	output	[11:0]  taps108x;
	output	[11:0]  taps109x;
	output	[11:0]  taps10x;
	output	[11:0]  taps110x;
	output	[11:0]  taps111x;
	output	[11:0]  taps112x;
	output	[11:0]  taps113x;
	output	[11:0]  taps114x;
	output	[11:0]  taps115x;
	output	[11:0]  taps116x;
	output	[11:0]  taps117x;
	output	[11:0]  taps118x;
	output	[11:0]  taps119x;
	output	[11:0]  taps11x;
	output	[11:0]  taps120x;
	output	[11:0]  taps121x;
	output	[11:0]  taps122x;
	output	[11:0]  taps123x;
	output	[11:0]  taps124x;
	output	[11:0]  taps125x;
	output	[11:0]  taps126x;
	output	[11:0]  taps127x;
	output	[11:0]  taps12x;
	output	[11:0]  taps13x;
	output	[11:0]  taps14x;
	output	[11:0]  taps15x;
	output	[11:0]  taps16x;
	output	[11:0]  taps17x;
	output	[11:0]  taps18x;
	output	[11:0]  taps19x;
	output	[11:0]  taps1x;
	output	[11:0]  taps20x;
	output	[11:0]  taps21x;
	output	[11:0]  taps22x;
	output	[11:0]  taps23x;
	output	[11:0]  taps24x;
	output	[11:0]  taps25x;
	output	[11:0]  taps26x;
	output	[11:0]  taps27x;
	output	[11:0]  taps28x;
	output	[11:0]  taps29x;
	output	[11:0]  taps2x;
	output	[11:0]  taps30x;
	output	[11:0]  taps31x;
	output	[11:0]  taps32x;
	output	[11:0]  taps33x;
	output	[11:0]  taps34x;
	output	[11:0]  taps35x;
	output	[11:0]  taps36x;
	output	[11:0]  taps37x;
	output	[11:0]  taps38x;
	output	[11:0]  taps39x;
	output	[11:0]  taps3x;
	output	[11:0]  taps40x;
	output	[11:0]  taps41x;
	output	[11:0]  taps42x;
	output	[11:0]  taps43x;
	output	[11:0]  taps44x;
	output	[11:0]  taps45x;
	output	[11:0]  taps46x;
	output	[11:0]  taps47x;
	output	[11:0]  taps48x;
	output	[11:0]  taps49x;
	output	[11:0]  taps4x;
	output	[11:0]  taps50x;
	output	[11:0]  taps51x;
	output	[11:0]  taps52x;
	output	[11:0]  taps53x;
	output	[11:0]  taps54x;
	output	[11:0]  taps55x;
	output	[11:0]  taps56x;
	output	[11:0]  taps57x;
	output	[11:0]  taps58x;
	output	[11:0]  taps59x;
	output	[11:0]  taps5x;
	output	[11:0]  taps60x;
	output	[11:0]  taps61x;
	output	[11:0]  taps62x;
	output	[11:0]  taps63x;
	output	[11:0]  taps64x;
	output	[11:0]  taps65x;
	output	[11:0]  taps66x;
	output	[11:0]  taps67x;
	output	[11:0]  taps68x;
	output	[11:0]  taps69x;
	output	[11:0]  taps6x;
	output	[11:0]  taps70x;
	output	[11:0]  taps71x;
	output	[11:0]  taps72x;
	output	[11:0]  taps73x;
	output	[11:0]  taps74x;
	output	[11:0]  taps75x;
	output	[11:0]  taps76x;
	output	[11:0]  taps77x;
	output	[11:0]  taps78x;
	output	[11:0]  taps79x;
	output	[11:0]  taps7x;
	output	[11:0]  taps80x;
	output	[11:0]  taps81x;
	output	[11:0]  taps82x;
	output	[11:0]  taps83x;
	output	[11:0]  taps84x;
	output	[11:0]  taps85x;
	output	[11:0]  taps86x;
	output	[11:0]  taps87x;
	output	[11:0]  taps88x;
	output	[11:0]  taps89x;
	output	[11:0]  taps8x;
	output	[11:0]  taps90x;
	output	[11:0]  taps91x;
	output	[11:0]  taps92x;
	output	[11:0]  taps93x;
	output	[11:0]  taps94x;
	output	[11:0]  taps95x;
	output	[11:0]  taps96x;
	output	[11:0]  taps97x;
	output	[11:0]  taps98x;
	output	[11:0]  taps99x;
	output	[11:0]  taps9x;

	wire [1535:0] sub_wire0;
	wire [11:0] sub_wire31;
	wire [1163:1152] sub_wire255 = sub_wire0[1163:1152];
	wire [947:936] sub_wire254 = sub_wire0[947:936];
	wire [947:936] sub_wire253 = sub_wire254[947:936];
	wire [1043:1032] sub_wire252 = sub_wire0[1043:1032];
	wire [1043:1032] sub_wire251 = sub_wire252[1043:1032];
	wire [827:816] sub_wire250 = sub_wire0[827:816];
	wire [827:816] sub_wire249 = sub_wire250[827:816];
	wire [1139:1128] sub_wire248 = sub_wire0[1139:1128];
	wire [1139:1128] sub_wire247 = sub_wire248[1139:1128];
	wire [923:912] sub_wire246 = sub_wire0[923:912];
	wire [923:912] sub_wire245 = sub_wire246[923:912];
	wire [707:696] sub_wire244 = sub_wire0[707:696];
	wire [707:696] sub_wire243 = sub_wire244[707:696];
	wire [1019:1008] sub_wire242 = sub_wire0[1019:1008];
	wire [1019:1008] sub_wire241 = sub_wire242[1019:1008];
	wire [803:792] sub_wire240 = sub_wire0[803:792];
	wire [803:792] sub_wire239 = sub_wire240[803:792];
	wire [587:576] sub_wire238 = sub_wire0[587:576];
	wire [587:576] sub_wire237 = sub_wire238[587:576];
	wire [1115:1104] sub_wire236 = sub_wire0[1115:1104];
	wire [1115:1104] sub_wire235 = sub_wire236[1115:1104];
	wire [899:888] sub_wire234 = sub_wire0[899:888];
	wire [899:888] sub_wire233 = sub_wire234[899:888];
	wire [683:672] sub_wire232 = sub_wire0[683:672];
	wire [683:672] sub_wire231 = sub_wire232[683:672];
	wire [467:456] sub_wire230 = sub_wire0[467:456];
	wire [467:456] sub_wire229 = sub_wire230[467:456];
	wire [995:984] sub_wire228 = sub_wire0[995:984];
	wire [995:984] sub_wire227 = sub_wire228[995:984];
	wire [779:768] sub_wire226 = sub_wire0[779:768];
	wire [779:768] sub_wire225 = sub_wire226[779:768];
	wire [563:552] sub_wire224 = sub_wire0[563:552];
	wire [563:552] sub_wire223 = sub_wire224[563:552];
	wire [347:336] sub_wire222 = sub_wire0[347:336];
	wire [347:336] sub_wire221 = sub_wire222[347:336];
	wire [1427:1416] sub_wire220 = sub_wire0[1427:1416];
	wire [1427:1416] sub_wire219 = sub_wire220[1427:1416];
	wire [119:108] sub_wire218 = sub_wire0[119:108];
	wire [119:108] sub_wire217 = sub_wire218[119:108];
	wire [1091:1080] sub_wire216 = sub_wire0[1091:1080];
	wire [1091:1080] sub_wire215 = sub_wire216[1091:1080];
	wire [875:864] sub_wire214 = sub_wire0[875:864];
	wire [875:864] sub_wire213 = sub_wire214[875:864];
	wire [659:648] sub_wire212 = sub_wire0[659:648];
	wire [659:648] sub_wire211 = sub_wire212[659:648];
	wire [443:432] sub_wire210 = sub_wire0[443:432];
	wire [443:432] sub_wire209 = sub_wire210[443:432];
	wire [227:216] sub_wire208 = sub_wire0[227:216];
	wire [227:216] sub_wire207 = sub_wire208[227:216];
	wire [1523:1512] sub_wire206 = sub_wire0[1523:1512];
	wire [1523:1512] sub_wire205 = sub_wire206[1523:1512];
	wire [1307:1296] sub_wire204 = sub_wire0[1307:1296];
	wire [1307:1296] sub_wire203 = sub_wire204[1307:1296];
	wire [971:960] sub_wire202 = sub_wire0[971:960];
	wire [971:960] sub_wire201 = sub_wire202[971:960];
	wire [755:744] sub_wire200 = sub_wire0[755:744];
	wire [755:744] sub_wire199 = sub_wire200[755:744];
	wire [539:528] sub_wire198 = sub_wire0[539:528];
	wire [539:528] sub_wire197 = sub_wire198[539:528];
	wire [323:312] sub_wire196 = sub_wire0[323:312];
	wire [323:312] sub_wire195 = sub_wire196[323:312];
	wire [1403:1392] sub_wire194 = sub_wire0[1403:1392];
	wire [1403:1392] sub_wire193 = sub_wire194[1403:1392];
	wire [95:84] sub_wire192 = sub_wire0[95:84];
	wire [95:84] sub_wire191 = sub_wire192[95:84];
	wire [851:840] sub_wire190 = sub_wire0[851:840];
	wire [851:840] sub_wire189 = sub_wire190[851:840];
	wire [635:624] sub_wire188 = sub_wire0[635:624];
	wire [635:624] sub_wire187 = sub_wire188[635:624];
	wire [419:408] sub_wire186 = sub_wire0[419:408];
	wire [419:408] sub_wire185 = sub_wire186[419:408];
	wire [203:192] sub_wire184 = sub_wire0[203:192];
	wire [203:192] sub_wire183 = sub_wire184[203:192];
	wire [1499:1488] sub_wire182 = sub_wire0[1499:1488];
	wire [1499:1488] sub_wire181 = sub_wire182[1499:1488];
	wire [1283:1272] sub_wire180 = sub_wire0[1283:1272];
	wire [1283:1272] sub_wire179 = sub_wire180[1283:1272];
	wire [731:720] sub_wire178 = sub_wire0[731:720];
	wire [731:720] sub_wire177 = sub_wire178[731:720];
	wire [515:504] sub_wire176 = sub_wire0[515:504];
	wire [515:504] sub_wire175 = sub_wire176[515:504];
	wire [299:288] sub_wire174 = sub_wire0[299:288];
	wire [299:288] sub_wire173 = sub_wire174[299:288];
	wire [1379:1368] sub_wire172 = sub_wire0[1379:1368];
	wire [1379:1368] sub_wire171 = sub_wire172[1379:1368];
	wire [71:60] sub_wire170 = sub_wire0[71:60];
	wire [71:60] sub_wire169 = sub_wire170[71:60];
	wire [611:600] sub_wire168 = sub_wire0[611:600];
	wire [611:600] sub_wire167 = sub_wire168[611:600];
	wire [395:384] sub_wire166 = sub_wire0[395:384];
	wire [395:384] sub_wire165 = sub_wire166[395:384];
	wire [179:168] sub_wire164 = sub_wire0[179:168];
	wire [179:168] sub_wire163 = sub_wire164[179:168];
	wire [1475:1464] sub_wire162 = sub_wire0[1475:1464];
	wire [1475:1464] sub_wire161 = sub_wire162[1475:1464];
	wire [1259:1248] sub_wire160 = sub_wire0[1259:1248];
	wire [1259:1248] sub_wire159 = sub_wire160[1259:1248];
	wire [491:480] sub_wire158 = sub_wire0[491:480];
	wire [491:480] sub_wire157 = sub_wire158[491:480];
	wire [275:264] sub_wire156 = sub_wire0[275:264];
	wire [275:264] sub_wire155 = sub_wire156[275:264];
	wire [1355:1344] sub_wire154 = sub_wire0[1355:1344];
	wire [1355:1344] sub_wire153 = sub_wire154[1355:1344];
	wire [47:36] sub_wire152 = sub_wire0[47:36];
	wire [47:36] sub_wire151 = sub_wire152[47:36];
	wire [371:360] sub_wire150 = sub_wire0[371:360];
	wire [371:360] sub_wire149 = sub_wire150[371:360];
	wire [155:144] sub_wire148 = sub_wire0[155:144];
	wire [155:144] sub_wire147 = sub_wire148[155:144];
	wire [1451:1440] sub_wire146 = sub_wire0[1451:1440];
	wire [1451:1440] sub_wire145 = sub_wire146[1451:1440];
	wire [1235:1224] sub_wire144 = sub_wire0[1235:1224];
	wire [1235:1224] sub_wire143 = sub_wire144[1235:1224];
	wire [1199:1188] sub_wire142 = sub_wire0[1199:1188];
	wire [1199:1188] sub_wire141 = sub_wire142[1199:1188];
	wire [251:240] sub_wire140 = sub_wire0[251:240];
	wire [251:240] sub_wire139 = sub_wire140[251:240];
	wire [1331:1320] sub_wire138 = sub_wire0[1331:1320];
	wire [1331:1320] sub_wire137 = sub_wire138[1331:1320];
	wire [1079:1068] sub_wire136 = sub_wire0[1079:1068];
	wire [1079:1068] sub_wire135 = sub_wire136[1079:1068];
	wire [23:12] sub_wire134 = sub_wire0[23:12];
	wire [23:12] sub_wire133 = sub_wire134[23:12];
	wire [131:120] sub_wire132 = sub_wire0[131:120];
	wire [131:120] sub_wire131 = sub_wire132[131:120];
	wire [1211:1200] sub_wire130 = sub_wire0[1211:1200];
	wire [1211:1200] sub_wire129 = sub_wire130[1211:1200];
	wire [1175:1164] sub_wire128 = sub_wire0[1175:1164];
	wire [1175:1164] sub_wire127 = sub_wire128[1175:1164];
	wire [959:948] sub_wire126 = sub_wire0[959:948];
	wire [959:948] sub_wire125 = sub_wire126[959:948];
	wire [1055:1044] sub_wire124 = sub_wire0[1055:1044];
	wire [1055:1044] sub_wire123 = sub_wire124[1055:1044];
	wire [839:828] sub_wire122 = sub_wire0[839:828];
	wire [839:828] sub_wire121 = sub_wire122[839:828];
	wire [1151:1140] sub_wire120 = sub_wire0[1151:1140];
	wire [1151:1140] sub_wire119 = sub_wire120[1151:1140];
	wire [935:924] sub_wire118 = sub_wire0[935:924];
	wire [935:924] sub_wire117 = sub_wire118[935:924];
	wire [719:708] sub_wire116 = sub_wire0[719:708];
	wire [719:708] sub_wire115 = sub_wire116[719:708];
	wire [1031:1020] sub_wire114 = sub_wire0[1031:1020];
	wire [1031:1020] sub_wire113 = sub_wire114[1031:1020];
	wire [815:804] sub_wire112 = sub_wire0[815:804];
	wire [815:804] sub_wire111 = sub_wire112[815:804];
	wire [599:588] sub_wire110 = sub_wire0[599:588];
	wire [599:588] sub_wire109 = sub_wire110[599:588];
	wire [1127:1116] sub_wire108 = sub_wire0[1127:1116];
	wire [1127:1116] sub_wire107 = sub_wire108[1127:1116];
	wire [911:900] sub_wire106 = sub_wire0[911:900];
	wire [911:900] sub_wire105 = sub_wire106[911:900];
	wire [695:684] sub_wire104 = sub_wire0[695:684];
	wire [695:684] sub_wire103 = sub_wire104[695:684];
	wire [479:468] sub_wire102 = sub_wire0[479:468];
	wire [479:468] sub_wire101 = sub_wire102[479:468];
	wire [1007:996] sub_wire100 = sub_wire0[1007:996];
	wire [1007:996] sub_wire99 = sub_wire100[1007:996];
	wire [791:780] sub_wire98 = sub_wire0[791:780];
	wire [791:780] sub_wire97 = sub_wire98[791:780];
	wire [575:564] sub_wire96 = sub_wire0[575:564];
	wire [575:564] sub_wire95 = sub_wire96[575:564];
	wire [359:348] sub_wire94 = sub_wire0[359:348];
	wire [359:348] sub_wire93 = sub_wire94[359:348];
	wire [1439:1428] sub_wire92 = sub_wire0[1439:1428];
	wire [1439:1428] sub_wire91 = sub_wire92[1439:1428];
	wire [1103:1092] sub_wire90 = sub_wire0[1103:1092];
	wire [1103:1092] sub_wire89 = sub_wire90[1103:1092];
	wire [887:876] sub_wire88 = sub_wire0[887:876];
	wire [887:876] sub_wire87 = sub_wire88[887:876];
	wire [671:660] sub_wire86 = sub_wire0[671:660];
	wire [671:660] sub_wire85 = sub_wire86[671:660];
	wire [455:444] sub_wire84 = sub_wire0[455:444];
	wire [455:444] sub_wire83 = sub_wire84[455:444];
	wire [239:228] sub_wire82 = sub_wire0[239:228];
	wire [239:228] sub_wire81 = sub_wire82[239:228];
	wire [1535:1524] sub_wire80 = sub_wire0[1535:1524];
	wire [1535:1524] sub_wire79 = sub_wire80[1535:1524];
	wire [1319:1308] sub_wire78 = sub_wire0[1319:1308];
	wire [1319:1308] sub_wire77 = sub_wire78[1319:1308];
	wire [983:972] sub_wire76 = sub_wire0[983:972];
	wire [983:972] sub_wire75 = sub_wire76[983:972];
	wire [767:756] sub_wire74 = sub_wire0[767:756];
	wire [767:756] sub_wire73 = sub_wire74[767:756];
	wire [551:540] sub_wire72 = sub_wire0[551:540];
	wire [551:540] sub_wire71 = sub_wire72[551:540];
	wire [335:324] sub_wire70 = sub_wire0[335:324];
	wire [335:324] sub_wire69 = sub_wire70[335:324];
	wire [1415:1404] sub_wire68 = sub_wire0[1415:1404];
	wire [1415:1404] sub_wire67 = sub_wire68[1415:1404];
	wire [107:96] sub_wire66 = sub_wire0[107:96];
	wire [107:96] sub_wire65 = sub_wire66[107:96];
	wire [863:852] sub_wire64 = sub_wire0[863:852];
	wire [863:852] sub_wire63 = sub_wire64[863:852];
	wire [647:636] sub_wire62 = sub_wire0[647:636];
	wire [647:636] sub_wire61 = sub_wire62[647:636];
	wire [431:420] sub_wire60 = sub_wire0[431:420];
	wire [431:420] sub_wire59 = sub_wire60[431:420];
	wire [215:204] sub_wire58 = sub_wire0[215:204];
	wire [215:204] sub_wire57 = sub_wire58[215:204];
	wire [1511:1500] sub_wire56 = sub_wire0[1511:1500];
	wire [1511:1500] sub_wire55 = sub_wire56[1511:1500];
	wire [1295:1284] sub_wire54 = sub_wire0[1295:1284];
	wire [1295:1284] sub_wire53 = sub_wire54[1295:1284];
	wire [743:732] sub_wire52 = sub_wire0[743:732];
	wire [743:732] sub_wire51 = sub_wire52[743:732];
	wire [527:516] sub_wire50 = sub_wire0[527:516];
	wire [527:516] sub_wire49 = sub_wire50[527:516];
	wire [311:300] sub_wire48 = sub_wire0[311:300];
	wire [311:300] sub_wire47 = sub_wire48[311:300];
	wire [1391:1380] sub_wire46 = sub_wire0[1391:1380];
	wire [1391:1380] sub_wire45 = sub_wire46[1391:1380];
	wire [83:72] sub_wire44 = sub_wire0[83:72];
	wire [83:72] sub_wire43 = sub_wire44[83:72];
	wire [623:612] sub_wire42 = sub_wire0[623:612];
	wire [623:612] sub_wire41 = sub_wire42[623:612];
	wire [407:396] sub_wire40 = sub_wire0[407:396];
	wire [407:396] sub_wire39 = sub_wire40[407:396];
	wire [191:180] sub_wire38 = sub_wire0[191:180];
	wire [191:180] sub_wire37 = sub_wire38[191:180];
	wire [1487:1476] sub_wire36 = sub_wire0[1487:1476];
	wire [1487:1476] sub_wire35 = sub_wire36[1487:1476];
	wire [1271:1260] sub_wire34 = sub_wire0[1271:1260];
	wire [1271:1260] sub_wire33 = sub_wire34[1271:1260];
	wire [503:492] sub_wire32 = sub_wire0[503:492];
	wire [503:492] sub_wire30 = sub_wire32[503:492];
	wire [287:276] sub_wire29 = sub_wire0[287:276];
	wire [287:276] sub_wire28 = sub_wire29[287:276];
	wire [1367:1356] sub_wire27 = sub_wire0[1367:1356];
	wire [1367:1356] sub_wire26 = sub_wire27[1367:1356];
	wire [59:48] sub_wire25 = sub_wire0[59:48];
	wire [59:48] sub_wire24 = sub_wire25[59:48];
	wire [383:372] sub_wire23 = sub_wire0[383:372];
	wire [383:372] sub_wire22 = sub_wire23[383:372];
	wire [167:156] sub_wire21 = sub_wire0[167:156];
	wire [167:156] sub_wire20 = sub_wire21[167:156];
	wire [1463:1452] sub_wire19 = sub_wire0[1463:1452];
	wire [1463:1452] sub_wire18 = sub_wire19[1463:1452];
	wire [1247:1236] sub_wire17 = sub_wire0[1247:1236];
	wire [1247:1236] sub_wire16 = sub_wire17[1247:1236];
	wire [263:252] sub_wire15 = sub_wire0[263:252];
	wire [263:252] sub_wire14 = sub_wire15[263:252];
	wire [1343:1332] sub_wire13 = sub_wire0[1343:1332];
	wire [1343:1332] sub_wire12 = sub_wire13[1343:1332];
	wire [35:24] sub_wire11 = sub_wire0[35:24];
	wire [35:24] sub_wire10 = sub_wire11[35:24];
	wire [143:132] sub_wire9 = sub_wire0[143:132];
	wire [143:132] sub_wire8 = sub_wire9[143:132];
	wire [1223:1212] sub_wire7 = sub_wire0[1223:1212];
	wire [1223:1212] sub_wire6 = sub_wire7[1223:1212];
	wire [1187:1176] sub_wire5 = sub_wire0[1187:1176];
	wire [1187:1176] sub_wire4 = sub_wire5[1187:1176];
	wire [1067:1056] sub_wire3 = sub_wire0[1067:1056];
	wire [1067:1056] sub_wire2 = sub_wire3[1067:1056];
	wire [11:0] sub_wire1 = sub_wire0[11:0];
	wire [11:0] taps0x = sub_wire1[11:0];
	wire [11:0] taps88x = sub_wire2[1067:1056];
	wire [11:0] taps98x = sub_wire4[1187:1176];
	wire [11:0] taps101x = sub_wire6[1223:1212];
	wire [11:0] taps11x = sub_wire8[143:132];
	wire [11:0] taps2x = sub_wire10[35:24];
	wire [11:0] taps111x = sub_wire12[1343:1332];
	wire [11:0] taps21x = sub_wire14[263:252];
	wire [11:0] taps103x = sub_wire16[1247:1236];
	wire [11:0] taps121x = sub_wire18[1463:1452];
	wire [11:0] taps13x = sub_wire20[167:156];
	wire [11:0] taps31x = sub_wire22[383:372];
	wire [11:0] taps4x = sub_wire24[59:48];
	wire [11:0] taps113x = sub_wire26[1367:1356];
	wire [11:0] taps23x = sub_wire28[287:276];
	wire [11:0] taps41x = sub_wire30[503:492];
	wire [11:0] shiftout = sub_wire31[11:0];
	wire [11:0] taps105x = sub_wire33[1271:1260];
	wire [11:0] taps123x = sub_wire35[1487:1476];
	wire [11:0] taps15x = sub_wire37[191:180];
	wire [11:0] taps33x = sub_wire39[407:396];
	wire [11:0] taps51x = sub_wire41[623:612];
	wire [11:0] taps6x = sub_wire43[83:72];
	wire [11:0] taps115x = sub_wire45[1391:1380];
	wire [11:0] taps25x = sub_wire47[311:300];
	wire [11:0] taps43x = sub_wire49[527:516];
	wire [11:0] taps61x = sub_wire51[743:732];
	wire [11:0] taps107x = sub_wire53[1295:1284];
	wire [11:0] taps125x = sub_wire55[1511:1500];
	wire [11:0] taps17x = sub_wire57[215:204];
	wire [11:0] taps35x = sub_wire59[431:420];
	wire [11:0] taps53x = sub_wire61[647:636];
	wire [11:0] taps71x = sub_wire63[863:852];
	wire [11:0] taps8x = sub_wire65[107:96];
	wire [11:0] taps117x = sub_wire67[1415:1404];
	wire [11:0] taps27x = sub_wire69[335:324];
	wire [11:0] taps45x = sub_wire71[551:540];
	wire [11:0] taps63x = sub_wire73[767:756];
	wire [11:0] taps81x = sub_wire75[983:972];
	wire [11:0] taps109x = sub_wire77[1319:1308];
	wire [11:0] taps127x = sub_wire79[1535:1524];
	wire [11:0] taps19x = sub_wire81[239:228];
	wire [11:0] taps37x = sub_wire83[455:444];
	wire [11:0] taps55x = sub_wire85[671:660];
	wire [11:0] taps73x = sub_wire87[887:876];
	wire [11:0] taps91x = sub_wire89[1103:1092];
	wire [11:0] taps119x = sub_wire91[1439:1428];
	wire [11:0] taps29x = sub_wire93[359:348];
	wire [11:0] taps47x = sub_wire95[575:564];
	wire [11:0] taps65x = sub_wire97[791:780];
	wire [11:0] taps83x = sub_wire99[1007:996];
	wire [11:0] taps39x = sub_wire101[479:468];
	wire [11:0] taps57x = sub_wire103[695:684];
	wire [11:0] taps75x = sub_wire105[911:900];
	wire [11:0] taps93x = sub_wire107[1127:1116];
	wire [11:0] taps49x = sub_wire109[599:588];
	wire [11:0] taps67x = sub_wire111[815:804];
	wire [11:0] taps85x = sub_wire113[1031:1020];
	wire [11:0] taps59x = sub_wire115[719:708];
	wire [11:0] taps77x = sub_wire117[935:924];
	wire [11:0] taps95x = sub_wire119[1151:1140];
	wire [11:0] taps69x = sub_wire121[839:828];
	wire [11:0] taps87x = sub_wire123[1055:1044];
	wire [11:0] taps79x = sub_wire125[959:948];
	wire [11:0] taps97x = sub_wire127[1175:1164];
	wire [11:0] taps100x = sub_wire129[1211:1200];
	wire [11:0] taps10x = sub_wire131[131:120];
	wire [11:0] taps1x = sub_wire133[23:12];
	wire [11:0] taps89x = sub_wire135[1079:1068];
	wire [11:0] taps110x = sub_wire137[1331:1320];
	wire [11:0] taps20x = sub_wire139[251:240];
	wire [11:0] taps99x = sub_wire141[1199:1188];
	wire [11:0] taps102x = sub_wire143[1235:1224];
	wire [11:0] taps120x = sub_wire145[1451:1440];
	wire [11:0] taps12x = sub_wire147[155:144];
	wire [11:0] taps30x = sub_wire149[371:360];
	wire [11:0] taps3x = sub_wire151[47:36];
	wire [11:0] taps112x = sub_wire153[1355:1344];
	wire [11:0] taps22x = sub_wire155[275:264];
	wire [11:0] taps40x = sub_wire157[491:480];
	wire [11:0] taps104x = sub_wire159[1259:1248];
	wire [11:0] taps122x = sub_wire161[1475:1464];
	wire [11:0] taps14x = sub_wire163[179:168];
	wire [11:0] taps32x = sub_wire165[395:384];
	wire [11:0] taps50x = sub_wire167[611:600];
	wire [11:0] taps5x = sub_wire169[71:60];
	wire [11:0] taps114x = sub_wire171[1379:1368];
	wire [11:0] taps24x = sub_wire173[299:288];
	wire [11:0] taps42x = sub_wire175[515:504];
	wire [11:0] taps60x = sub_wire177[731:720];
	wire [11:0] taps106x = sub_wire179[1283:1272];
	wire [11:0] taps124x = sub_wire181[1499:1488];
	wire [11:0] taps16x = sub_wire183[203:192];
	wire [11:0] taps34x = sub_wire185[419:408];
	wire [11:0] taps52x = sub_wire187[635:624];
	wire [11:0] taps70x = sub_wire189[851:840];
	wire [11:0] taps7x = sub_wire191[95:84];
	wire [11:0] taps116x = sub_wire193[1403:1392];
	wire [11:0] taps26x = sub_wire195[323:312];
	wire [11:0] taps44x = sub_wire197[539:528];
	wire [11:0] taps62x = sub_wire199[755:744];
	wire [11:0] taps80x = sub_wire201[971:960];
	wire [11:0] taps108x = sub_wire203[1307:1296];
	wire [11:0] taps126x = sub_wire205[1523:1512];
	wire [11:0] taps18x = sub_wire207[227:216];
	wire [11:0] taps36x = sub_wire209[443:432];
	wire [11:0] taps54x = sub_wire211[659:648];
	wire [11:0] taps72x = sub_wire213[875:864];
	wire [11:0] taps90x = sub_wire215[1091:1080];
	wire [11:0] taps9x = sub_wire217[119:108];
	wire [11:0] taps118x = sub_wire219[1427:1416];
	wire [11:0] taps28x = sub_wire221[347:336];
	wire [11:0] taps46x = sub_wire223[563:552];
	wire [11:0] taps64x = sub_wire225[779:768];
	wire [11:0] taps82x = sub_wire227[995:984];
	wire [11:0] taps38x = sub_wire229[467:456];
	wire [11:0] taps56x = sub_wire231[683:672];
	wire [11:0] taps74x = sub_wire233[899:888];
	wire [11:0] taps92x = sub_wire235[1115:1104];
	wire [11:0] taps48x = sub_wire237[587:576];
	wire [11:0] taps66x = sub_wire239[803:792];
	wire [11:0] taps84x = sub_wire241[1019:1008];
	wire [11:0] taps58x = sub_wire243[707:696];
	wire [11:0] taps76x = sub_wire245[923:912];
	wire [11:0] taps94x = sub_wire247[1139:1128];
	wire [11:0] taps68x = sub_wire249[827:816];
	wire [11:0] taps86x = sub_wire251[1043:1032];
	wire [11:0] taps78x = sub_wire253[947:936];
	wire [11:0] taps96x = sub_wire255[1163:1152];

	altshift_taps	ALTSHIFT_TAPS_component (
				.clock (clock),
				.shiftin (shiftin),
				.taps (sub_wire0),
				.shiftout (sub_wire31)
				// synopsys translate_off
				,
				.aclr (),
				.clken ()
				// synopsys translate_on
				);
	defparam
		ALTSHIFT_TAPS_component.intended_device_family = "Cyclone IV E",
		ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=AUTO",
		ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
		ALTSHIFT_TAPS_component.number_of_taps = 128,
		ALTSHIFT_TAPS_component.tap_distance = 3,
		ALTSHIFT_TAPS_component.width = 12;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "0"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "128"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "3"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "3"
// Retrieval info: PRIVATE: WIDTH NUMERIC "12"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=AUTO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "128"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "3"
// Retrieval info: CONSTANT: WIDTH NUMERIC "12"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 12 0 INPUT NODEFVAL "shiftin[11..0]"
// Retrieval info: USED_PORT: shiftout 0 0 12 0 OUTPUT NODEFVAL "shiftout[11..0]"
// Retrieval info: USED_PORT: taps0x 0 0 12 0 OUTPUT NODEFVAL "taps0x[11..0]"
// Retrieval info: USED_PORT: taps100x 0 0 12 0 OUTPUT NODEFVAL "taps100x[11..0]"
// Retrieval info: USED_PORT: taps101x 0 0 12 0 OUTPUT NODEFVAL "taps101x[11..0]"
// Retrieval info: USED_PORT: taps102x 0 0 12 0 OUTPUT NODEFVAL "taps102x[11..0]"
// Retrieval info: USED_PORT: taps103x 0 0 12 0 OUTPUT NODEFVAL "taps103x[11..0]"
// Retrieval info: USED_PORT: taps104x 0 0 12 0 OUTPUT NODEFVAL "taps104x[11..0]"
// Retrieval info: USED_PORT: taps105x 0 0 12 0 OUTPUT NODEFVAL "taps105x[11..0]"
// Retrieval info: USED_PORT: taps106x 0 0 12 0 OUTPUT NODEFVAL "taps106x[11..0]"
// Retrieval info: USED_PORT: taps107x 0 0 12 0 OUTPUT NODEFVAL "taps107x[11..0]"
// Retrieval info: USED_PORT: taps108x 0 0 12 0 OUTPUT NODEFVAL "taps108x[11..0]"
// Retrieval info: USED_PORT: taps109x 0 0 12 0 OUTPUT NODEFVAL "taps109x[11..0]"
// Retrieval info: USED_PORT: taps10x 0 0 12 0 OUTPUT NODEFVAL "taps10x[11..0]"
// Retrieval info: USED_PORT: taps110x 0 0 12 0 OUTPUT NODEFVAL "taps110x[11..0]"
// Retrieval info: USED_PORT: taps111x 0 0 12 0 OUTPUT NODEFVAL "taps111x[11..0]"
// Retrieval info: USED_PORT: taps112x 0 0 12 0 OUTPUT NODEFVAL "taps112x[11..0]"
// Retrieval info: USED_PORT: taps113x 0 0 12 0 OUTPUT NODEFVAL "taps113x[11..0]"
// Retrieval info: USED_PORT: taps114x 0 0 12 0 OUTPUT NODEFVAL "taps114x[11..0]"
// Retrieval info: USED_PORT: taps115x 0 0 12 0 OUTPUT NODEFVAL "taps115x[11..0]"
// Retrieval info: USED_PORT: taps116x 0 0 12 0 OUTPUT NODEFVAL "taps116x[11..0]"
// Retrieval info: USED_PORT: taps117x 0 0 12 0 OUTPUT NODEFVAL "taps117x[11..0]"
// Retrieval info: USED_PORT: taps118x 0 0 12 0 OUTPUT NODEFVAL "taps118x[11..0]"
// Retrieval info: USED_PORT: taps119x 0 0 12 0 OUTPUT NODEFVAL "taps119x[11..0]"
// Retrieval info: USED_PORT: taps11x 0 0 12 0 OUTPUT NODEFVAL "taps11x[11..0]"
// Retrieval info: USED_PORT: taps120x 0 0 12 0 OUTPUT NODEFVAL "taps120x[11..0]"
// Retrieval info: USED_PORT: taps121x 0 0 12 0 OUTPUT NODEFVAL "taps121x[11..0]"
// Retrieval info: USED_PORT: taps122x 0 0 12 0 OUTPUT NODEFVAL "taps122x[11..0]"
// Retrieval info: USED_PORT: taps123x 0 0 12 0 OUTPUT NODEFVAL "taps123x[11..0]"
// Retrieval info: USED_PORT: taps124x 0 0 12 0 OUTPUT NODEFVAL "taps124x[11..0]"
// Retrieval info: USED_PORT: taps125x 0 0 12 0 OUTPUT NODEFVAL "taps125x[11..0]"
// Retrieval info: USED_PORT: taps126x 0 0 12 0 OUTPUT NODEFVAL "taps126x[11..0]"
// Retrieval info: USED_PORT: taps127x 0 0 12 0 OUTPUT NODEFVAL "taps127x[11..0]"
// Retrieval info: USED_PORT: taps12x 0 0 12 0 OUTPUT NODEFVAL "taps12x[11..0]"
// Retrieval info: USED_PORT: taps13x 0 0 12 0 OUTPUT NODEFVAL "taps13x[11..0]"
// Retrieval info: USED_PORT: taps14x 0 0 12 0 OUTPUT NODEFVAL "taps14x[11..0]"
// Retrieval info: USED_PORT: taps15x 0 0 12 0 OUTPUT NODEFVAL "taps15x[11..0]"
// Retrieval info: USED_PORT: taps16x 0 0 12 0 OUTPUT NODEFVAL "taps16x[11..0]"
// Retrieval info: USED_PORT: taps17x 0 0 12 0 OUTPUT NODEFVAL "taps17x[11..0]"
// Retrieval info: USED_PORT: taps18x 0 0 12 0 OUTPUT NODEFVAL "taps18x[11..0]"
// Retrieval info: USED_PORT: taps19x 0 0 12 0 OUTPUT NODEFVAL "taps19x[11..0]"
// Retrieval info: USED_PORT: taps1x 0 0 12 0 OUTPUT NODEFVAL "taps1x[11..0]"
// Retrieval info: USED_PORT: taps20x 0 0 12 0 OUTPUT NODEFVAL "taps20x[11..0]"
// Retrieval info: USED_PORT: taps21x 0 0 12 0 OUTPUT NODEFVAL "taps21x[11..0]"
// Retrieval info: USED_PORT: taps22x 0 0 12 0 OUTPUT NODEFVAL "taps22x[11..0]"
// Retrieval info: USED_PORT: taps23x 0 0 12 0 OUTPUT NODEFVAL "taps23x[11..0]"
// Retrieval info: USED_PORT: taps24x 0 0 12 0 OUTPUT NODEFVAL "taps24x[11..0]"
// Retrieval info: USED_PORT: taps25x 0 0 12 0 OUTPUT NODEFVAL "taps25x[11..0]"
// Retrieval info: USED_PORT: taps26x 0 0 12 0 OUTPUT NODEFVAL "taps26x[11..0]"
// Retrieval info: USED_PORT: taps27x 0 0 12 0 OUTPUT NODEFVAL "taps27x[11..0]"
// Retrieval info: USED_PORT: taps28x 0 0 12 0 OUTPUT NODEFVAL "taps28x[11..0]"
// Retrieval info: USED_PORT: taps29x 0 0 12 0 OUTPUT NODEFVAL "taps29x[11..0]"
// Retrieval info: USED_PORT: taps2x 0 0 12 0 OUTPUT NODEFVAL "taps2x[11..0]"
// Retrieval info: USED_PORT: taps30x 0 0 12 0 OUTPUT NODEFVAL "taps30x[11..0]"
// Retrieval info: USED_PORT: taps31x 0 0 12 0 OUTPUT NODEFVAL "taps31x[11..0]"
// Retrieval info: USED_PORT: taps32x 0 0 12 0 OUTPUT NODEFVAL "taps32x[11..0]"
// Retrieval info: USED_PORT: taps33x 0 0 12 0 OUTPUT NODEFVAL "taps33x[11..0]"
// Retrieval info: USED_PORT: taps34x 0 0 12 0 OUTPUT NODEFVAL "taps34x[11..0]"
// Retrieval info: USED_PORT: taps35x 0 0 12 0 OUTPUT NODEFVAL "taps35x[11..0]"
// Retrieval info: USED_PORT: taps36x 0 0 12 0 OUTPUT NODEFVAL "taps36x[11..0]"
// Retrieval info: USED_PORT: taps37x 0 0 12 0 OUTPUT NODEFVAL "taps37x[11..0]"
// Retrieval info: USED_PORT: taps38x 0 0 12 0 OUTPUT NODEFVAL "taps38x[11..0]"
// Retrieval info: USED_PORT: taps39x 0 0 12 0 OUTPUT NODEFVAL "taps39x[11..0]"
// Retrieval info: USED_PORT: taps3x 0 0 12 0 OUTPUT NODEFVAL "taps3x[11..0]"
// Retrieval info: USED_PORT: taps40x 0 0 12 0 OUTPUT NODEFVAL "taps40x[11..0]"
// Retrieval info: USED_PORT: taps41x 0 0 12 0 OUTPUT NODEFVAL "taps41x[11..0]"
// Retrieval info: USED_PORT: taps42x 0 0 12 0 OUTPUT NODEFVAL "taps42x[11..0]"
// Retrieval info: USED_PORT: taps43x 0 0 12 0 OUTPUT NODEFVAL "taps43x[11..0]"
// Retrieval info: USED_PORT: taps44x 0 0 12 0 OUTPUT NODEFVAL "taps44x[11..0]"
// Retrieval info: USED_PORT: taps45x 0 0 12 0 OUTPUT NODEFVAL "taps45x[11..0]"
// Retrieval info: USED_PORT: taps46x 0 0 12 0 OUTPUT NODEFVAL "taps46x[11..0]"
// Retrieval info: USED_PORT: taps47x 0 0 12 0 OUTPUT NODEFVAL "taps47x[11..0]"
// Retrieval info: USED_PORT: taps48x 0 0 12 0 OUTPUT NODEFVAL "taps48x[11..0]"
// Retrieval info: USED_PORT: taps49x 0 0 12 0 OUTPUT NODEFVAL "taps49x[11..0]"
// Retrieval info: USED_PORT: taps4x 0 0 12 0 OUTPUT NODEFVAL "taps4x[11..0]"
// Retrieval info: USED_PORT: taps50x 0 0 12 0 OUTPUT NODEFVAL "taps50x[11..0]"
// Retrieval info: USED_PORT: taps51x 0 0 12 0 OUTPUT NODEFVAL "taps51x[11..0]"
// Retrieval info: USED_PORT: taps52x 0 0 12 0 OUTPUT NODEFVAL "taps52x[11..0]"
// Retrieval info: USED_PORT: taps53x 0 0 12 0 OUTPUT NODEFVAL "taps53x[11..0]"
// Retrieval info: USED_PORT: taps54x 0 0 12 0 OUTPUT NODEFVAL "taps54x[11..0]"
// Retrieval info: USED_PORT: taps55x 0 0 12 0 OUTPUT NODEFVAL "taps55x[11..0]"
// Retrieval info: USED_PORT: taps56x 0 0 12 0 OUTPUT NODEFVAL "taps56x[11..0]"
// Retrieval info: USED_PORT: taps57x 0 0 12 0 OUTPUT NODEFVAL "taps57x[11..0]"
// Retrieval info: USED_PORT: taps58x 0 0 12 0 OUTPUT NODEFVAL "taps58x[11..0]"
// Retrieval info: USED_PORT: taps59x 0 0 12 0 OUTPUT NODEFVAL "taps59x[11..0]"
// Retrieval info: USED_PORT: taps5x 0 0 12 0 OUTPUT NODEFVAL "taps5x[11..0]"
// Retrieval info: USED_PORT: taps60x 0 0 12 0 OUTPUT NODEFVAL "taps60x[11..0]"
// Retrieval info: USED_PORT: taps61x 0 0 12 0 OUTPUT NODEFVAL "taps61x[11..0]"
// Retrieval info: USED_PORT: taps62x 0 0 12 0 OUTPUT NODEFVAL "taps62x[11..0]"
// Retrieval info: USED_PORT: taps63x 0 0 12 0 OUTPUT NODEFVAL "taps63x[11..0]"
// Retrieval info: USED_PORT: taps64x 0 0 12 0 OUTPUT NODEFVAL "taps64x[11..0]"
// Retrieval info: USED_PORT: taps65x 0 0 12 0 OUTPUT NODEFVAL "taps65x[11..0]"
// Retrieval info: USED_PORT: taps66x 0 0 12 0 OUTPUT NODEFVAL "taps66x[11..0]"
// Retrieval info: USED_PORT: taps67x 0 0 12 0 OUTPUT NODEFVAL "taps67x[11..0]"
// Retrieval info: USED_PORT: taps68x 0 0 12 0 OUTPUT NODEFVAL "taps68x[11..0]"
// Retrieval info: USED_PORT: taps69x 0 0 12 0 OUTPUT NODEFVAL "taps69x[11..0]"
// Retrieval info: USED_PORT: taps6x 0 0 12 0 OUTPUT NODEFVAL "taps6x[11..0]"
// Retrieval info: USED_PORT: taps70x 0 0 12 0 OUTPUT NODEFVAL "taps70x[11..0]"
// Retrieval info: USED_PORT: taps71x 0 0 12 0 OUTPUT NODEFVAL "taps71x[11..0]"
// Retrieval info: USED_PORT: taps72x 0 0 12 0 OUTPUT NODEFVAL "taps72x[11..0]"
// Retrieval info: USED_PORT: taps73x 0 0 12 0 OUTPUT NODEFVAL "taps73x[11..0]"
// Retrieval info: USED_PORT: taps74x 0 0 12 0 OUTPUT NODEFVAL "taps74x[11..0]"
// Retrieval info: USED_PORT: taps75x 0 0 12 0 OUTPUT NODEFVAL "taps75x[11..0]"
// Retrieval info: USED_PORT: taps76x 0 0 12 0 OUTPUT NODEFVAL "taps76x[11..0]"
// Retrieval info: USED_PORT: taps77x 0 0 12 0 OUTPUT NODEFVAL "taps77x[11..0]"
// Retrieval info: USED_PORT: taps78x 0 0 12 0 OUTPUT NODEFVAL "taps78x[11..0]"
// Retrieval info: USED_PORT: taps79x 0 0 12 0 OUTPUT NODEFVAL "taps79x[11..0]"
// Retrieval info: USED_PORT: taps7x 0 0 12 0 OUTPUT NODEFVAL "taps7x[11..0]"
// Retrieval info: USED_PORT: taps80x 0 0 12 0 OUTPUT NODEFVAL "taps80x[11..0]"
// Retrieval info: USED_PORT: taps81x 0 0 12 0 OUTPUT NODEFVAL "taps81x[11..0]"
// Retrieval info: USED_PORT: taps82x 0 0 12 0 OUTPUT NODEFVAL "taps82x[11..0]"
// Retrieval info: USED_PORT: taps83x 0 0 12 0 OUTPUT NODEFVAL "taps83x[11..0]"
// Retrieval info: USED_PORT: taps84x 0 0 12 0 OUTPUT NODEFVAL "taps84x[11..0]"
// Retrieval info: USED_PORT: taps85x 0 0 12 0 OUTPUT NODEFVAL "taps85x[11..0]"
// Retrieval info: USED_PORT: taps86x 0 0 12 0 OUTPUT NODEFVAL "taps86x[11..0]"
// Retrieval info: USED_PORT: taps87x 0 0 12 0 OUTPUT NODEFVAL "taps87x[11..0]"
// Retrieval info: USED_PORT: taps88x 0 0 12 0 OUTPUT NODEFVAL "taps88x[11..0]"
// Retrieval info: USED_PORT: taps89x 0 0 12 0 OUTPUT NODEFVAL "taps89x[11..0]"
// Retrieval info: USED_PORT: taps8x 0 0 12 0 OUTPUT NODEFVAL "taps8x[11..0]"
// Retrieval info: USED_PORT: taps90x 0 0 12 0 OUTPUT NODEFVAL "taps90x[11..0]"
// Retrieval info: USED_PORT: taps91x 0 0 12 0 OUTPUT NODEFVAL "taps91x[11..0]"
// Retrieval info: USED_PORT: taps92x 0 0 12 0 OUTPUT NODEFVAL "taps92x[11..0]"
// Retrieval info: USED_PORT: taps93x 0 0 12 0 OUTPUT NODEFVAL "taps93x[11..0]"
// Retrieval info: USED_PORT: taps94x 0 0 12 0 OUTPUT NODEFVAL "taps94x[11..0]"
// Retrieval info: USED_PORT: taps95x 0 0 12 0 OUTPUT NODEFVAL "taps95x[11..0]"
// Retrieval info: USED_PORT: taps96x 0 0 12 0 OUTPUT NODEFVAL "taps96x[11..0]"
// Retrieval info: USED_PORT: taps97x 0 0 12 0 OUTPUT NODEFVAL "taps97x[11..0]"
// Retrieval info: USED_PORT: taps98x 0 0 12 0 OUTPUT NODEFVAL "taps98x[11..0]"
// Retrieval info: USED_PORT: taps99x 0 0 12 0 OUTPUT NODEFVAL "taps99x[11..0]"
// Retrieval info: USED_PORT: taps9x 0 0 12 0 OUTPUT NODEFVAL "taps9x[11..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 12 0 shiftin 0 0 12 0
// Retrieval info: CONNECT: shiftout 0 0 12 0 @shiftout 0 0 12 0
// Retrieval info: CONNECT: taps0x 0 0 12 0 @taps 0 0 12 0
// Retrieval info: CONNECT: taps100x 0 0 12 0 @taps 0 0 12 1200
// Retrieval info: CONNECT: taps101x 0 0 12 0 @taps 0 0 12 1212
// Retrieval info: CONNECT: taps102x 0 0 12 0 @taps 0 0 12 1224
// Retrieval info: CONNECT: taps103x 0 0 12 0 @taps 0 0 12 1236
// Retrieval info: CONNECT: taps104x 0 0 12 0 @taps 0 0 12 1248
// Retrieval info: CONNECT: taps105x 0 0 12 0 @taps 0 0 12 1260
// Retrieval info: CONNECT: taps106x 0 0 12 0 @taps 0 0 12 1272
// Retrieval info: CONNECT: taps107x 0 0 12 0 @taps 0 0 12 1284
// Retrieval info: CONNECT: taps108x 0 0 12 0 @taps 0 0 12 1296
// Retrieval info: CONNECT: taps109x 0 0 12 0 @taps 0 0 12 1308
// Retrieval info: CONNECT: taps10x 0 0 12 0 @taps 0 0 12 120
// Retrieval info: CONNECT: taps110x 0 0 12 0 @taps 0 0 12 1320
// Retrieval info: CONNECT: taps111x 0 0 12 0 @taps 0 0 12 1332
// Retrieval info: CONNECT: taps112x 0 0 12 0 @taps 0 0 12 1344
// Retrieval info: CONNECT: taps113x 0 0 12 0 @taps 0 0 12 1356
// Retrieval info: CONNECT: taps114x 0 0 12 0 @taps 0 0 12 1368
// Retrieval info: CONNECT: taps115x 0 0 12 0 @taps 0 0 12 1380
// Retrieval info: CONNECT: taps116x 0 0 12 0 @taps 0 0 12 1392
// Retrieval info: CONNECT: taps117x 0 0 12 0 @taps 0 0 12 1404
// Retrieval info: CONNECT: taps118x 0 0 12 0 @taps 0 0 12 1416
// Retrieval info: CONNECT: taps119x 0 0 12 0 @taps 0 0 12 1428
// Retrieval info: CONNECT: taps11x 0 0 12 0 @taps 0 0 12 132
// Retrieval info: CONNECT: taps120x 0 0 12 0 @taps 0 0 12 1440
// Retrieval info: CONNECT: taps121x 0 0 12 0 @taps 0 0 12 1452
// Retrieval info: CONNECT: taps122x 0 0 12 0 @taps 0 0 12 1464
// Retrieval info: CONNECT: taps123x 0 0 12 0 @taps 0 0 12 1476
// Retrieval info: CONNECT: taps124x 0 0 12 0 @taps 0 0 12 1488
// Retrieval info: CONNECT: taps125x 0 0 12 0 @taps 0 0 12 1500
// Retrieval info: CONNECT: taps126x 0 0 12 0 @taps 0 0 12 1512
// Retrieval info: CONNECT: taps127x 0 0 12 0 @taps 0 0 12 1524
// Retrieval info: CONNECT: taps12x 0 0 12 0 @taps 0 0 12 144
// Retrieval info: CONNECT: taps13x 0 0 12 0 @taps 0 0 12 156
// Retrieval info: CONNECT: taps14x 0 0 12 0 @taps 0 0 12 168
// Retrieval info: CONNECT: taps15x 0 0 12 0 @taps 0 0 12 180
// Retrieval info: CONNECT: taps16x 0 0 12 0 @taps 0 0 12 192
// Retrieval info: CONNECT: taps17x 0 0 12 0 @taps 0 0 12 204
// Retrieval info: CONNECT: taps18x 0 0 12 0 @taps 0 0 12 216
// Retrieval info: CONNECT: taps19x 0 0 12 0 @taps 0 0 12 228
// Retrieval info: CONNECT: taps1x 0 0 12 0 @taps 0 0 12 12
// Retrieval info: CONNECT: taps20x 0 0 12 0 @taps 0 0 12 240
// Retrieval info: CONNECT: taps21x 0 0 12 0 @taps 0 0 12 252
// Retrieval info: CONNECT: taps22x 0 0 12 0 @taps 0 0 12 264
// Retrieval info: CONNECT: taps23x 0 0 12 0 @taps 0 0 12 276
// Retrieval info: CONNECT: taps24x 0 0 12 0 @taps 0 0 12 288
// Retrieval info: CONNECT: taps25x 0 0 12 0 @taps 0 0 12 300
// Retrieval info: CONNECT: taps26x 0 0 12 0 @taps 0 0 12 312
// Retrieval info: CONNECT: taps27x 0 0 12 0 @taps 0 0 12 324
// Retrieval info: CONNECT: taps28x 0 0 12 0 @taps 0 0 12 336
// Retrieval info: CONNECT: taps29x 0 0 12 0 @taps 0 0 12 348
// Retrieval info: CONNECT: taps2x 0 0 12 0 @taps 0 0 12 24
// Retrieval info: CONNECT: taps30x 0 0 12 0 @taps 0 0 12 360
// Retrieval info: CONNECT: taps31x 0 0 12 0 @taps 0 0 12 372
// Retrieval info: CONNECT: taps32x 0 0 12 0 @taps 0 0 12 384
// Retrieval info: CONNECT: taps33x 0 0 12 0 @taps 0 0 12 396
// Retrieval info: CONNECT: taps34x 0 0 12 0 @taps 0 0 12 408
// Retrieval info: CONNECT: taps35x 0 0 12 0 @taps 0 0 12 420
// Retrieval info: CONNECT: taps36x 0 0 12 0 @taps 0 0 12 432
// Retrieval info: CONNECT: taps37x 0 0 12 0 @taps 0 0 12 444
// Retrieval info: CONNECT: taps38x 0 0 12 0 @taps 0 0 12 456
// Retrieval info: CONNECT: taps39x 0 0 12 0 @taps 0 0 12 468
// Retrieval info: CONNECT: taps3x 0 0 12 0 @taps 0 0 12 36
// Retrieval info: CONNECT: taps40x 0 0 12 0 @taps 0 0 12 480
// Retrieval info: CONNECT: taps41x 0 0 12 0 @taps 0 0 12 492
// Retrieval info: CONNECT: taps42x 0 0 12 0 @taps 0 0 12 504
// Retrieval info: CONNECT: taps43x 0 0 12 0 @taps 0 0 12 516
// Retrieval info: CONNECT: taps44x 0 0 12 0 @taps 0 0 12 528
// Retrieval info: CONNECT: taps45x 0 0 12 0 @taps 0 0 12 540
// Retrieval info: CONNECT: taps46x 0 0 12 0 @taps 0 0 12 552
// Retrieval info: CONNECT: taps47x 0 0 12 0 @taps 0 0 12 564
// Retrieval info: CONNECT: taps48x 0 0 12 0 @taps 0 0 12 576
// Retrieval info: CONNECT: taps49x 0 0 12 0 @taps 0 0 12 588
// Retrieval info: CONNECT: taps4x 0 0 12 0 @taps 0 0 12 48
// Retrieval info: CONNECT: taps50x 0 0 12 0 @taps 0 0 12 600
// Retrieval info: CONNECT: taps51x 0 0 12 0 @taps 0 0 12 612
// Retrieval info: CONNECT: taps52x 0 0 12 0 @taps 0 0 12 624
// Retrieval info: CONNECT: taps53x 0 0 12 0 @taps 0 0 12 636
// Retrieval info: CONNECT: taps54x 0 0 12 0 @taps 0 0 12 648
// Retrieval info: CONNECT: taps55x 0 0 12 0 @taps 0 0 12 660
// Retrieval info: CONNECT: taps56x 0 0 12 0 @taps 0 0 12 672
// Retrieval info: CONNECT: taps57x 0 0 12 0 @taps 0 0 12 684
// Retrieval info: CONNECT: taps58x 0 0 12 0 @taps 0 0 12 696
// Retrieval info: CONNECT: taps59x 0 0 12 0 @taps 0 0 12 708
// Retrieval info: CONNECT: taps5x 0 0 12 0 @taps 0 0 12 60
// Retrieval info: CONNECT: taps60x 0 0 12 0 @taps 0 0 12 720
// Retrieval info: CONNECT: taps61x 0 0 12 0 @taps 0 0 12 732
// Retrieval info: CONNECT: taps62x 0 0 12 0 @taps 0 0 12 744
// Retrieval info: CONNECT: taps63x 0 0 12 0 @taps 0 0 12 756
// Retrieval info: CONNECT: taps64x 0 0 12 0 @taps 0 0 12 768
// Retrieval info: CONNECT: taps65x 0 0 12 0 @taps 0 0 12 780
// Retrieval info: CONNECT: taps66x 0 0 12 0 @taps 0 0 12 792
// Retrieval info: CONNECT: taps67x 0 0 12 0 @taps 0 0 12 804
// Retrieval info: CONNECT: taps68x 0 0 12 0 @taps 0 0 12 816
// Retrieval info: CONNECT: taps69x 0 0 12 0 @taps 0 0 12 828
// Retrieval info: CONNECT: taps6x 0 0 12 0 @taps 0 0 12 72
// Retrieval info: CONNECT: taps70x 0 0 12 0 @taps 0 0 12 840
// Retrieval info: CONNECT: taps71x 0 0 12 0 @taps 0 0 12 852
// Retrieval info: CONNECT: taps72x 0 0 12 0 @taps 0 0 12 864
// Retrieval info: CONNECT: taps73x 0 0 12 0 @taps 0 0 12 876
// Retrieval info: CONNECT: taps74x 0 0 12 0 @taps 0 0 12 888
// Retrieval info: CONNECT: taps75x 0 0 12 0 @taps 0 0 12 900
// Retrieval info: CONNECT: taps76x 0 0 12 0 @taps 0 0 12 912
// Retrieval info: CONNECT: taps77x 0 0 12 0 @taps 0 0 12 924
// Retrieval info: CONNECT: taps78x 0 0 12 0 @taps 0 0 12 936
// Retrieval info: CONNECT: taps79x 0 0 12 0 @taps 0 0 12 948
// Retrieval info: CONNECT: taps7x 0 0 12 0 @taps 0 0 12 84
// Retrieval info: CONNECT: taps80x 0 0 12 0 @taps 0 0 12 960
// Retrieval info: CONNECT: taps81x 0 0 12 0 @taps 0 0 12 972
// Retrieval info: CONNECT: taps82x 0 0 12 0 @taps 0 0 12 984
// Retrieval info: CONNECT: taps83x 0 0 12 0 @taps 0 0 12 996
// Retrieval info: CONNECT: taps84x 0 0 12 0 @taps 0 0 12 1008
// Retrieval info: CONNECT: taps85x 0 0 12 0 @taps 0 0 12 1020
// Retrieval info: CONNECT: taps86x 0 0 12 0 @taps 0 0 12 1032
// Retrieval info: CONNECT: taps87x 0 0 12 0 @taps 0 0 12 1044
// Retrieval info: CONNECT: taps88x 0 0 12 0 @taps 0 0 12 1056
// Retrieval info: CONNECT: taps89x 0 0 12 0 @taps 0 0 12 1068
// Retrieval info: CONNECT: taps8x 0 0 12 0 @taps 0 0 12 96
// Retrieval info: CONNECT: taps90x 0 0 12 0 @taps 0 0 12 1080
// Retrieval info: CONNECT: taps91x 0 0 12 0 @taps 0 0 12 1092
// Retrieval info: CONNECT: taps92x 0 0 12 0 @taps 0 0 12 1104
// Retrieval info: CONNECT: taps93x 0 0 12 0 @taps 0 0 12 1116
// Retrieval info: CONNECT: taps94x 0 0 12 0 @taps 0 0 12 1128
// Retrieval info: CONNECT: taps95x 0 0 12 0 @taps 0 0 12 1140
// Retrieval info: CONNECT: taps96x 0 0 12 0 @taps 0 0 12 1152
// Retrieval info: CONNECT: taps97x 0 0 12 0 @taps 0 0 12 1164
// Retrieval info: CONNECT: taps98x 0 0 12 0 @taps 0 0 12 1176
// Retrieval info: CONNECT: taps99x 0 0 12 0 @taps 0 0 12 1188
// Retrieval info: CONNECT: taps9x 0 0 12 0 @taps 0 0 12 108
// Retrieval info: GEN_FILE: TYPE_NORMAL history_reg.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL history_reg.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL history_reg.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL history_reg.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL history_reg_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL history_reg_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
